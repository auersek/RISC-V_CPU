`ifndef DEF_SV
`define DEF_SV

`define ALU_OPCODE_ADD =        4'b0000;
`define ALU_OPCODE_SUB =        4'b0001;

`endif
